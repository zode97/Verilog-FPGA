// TCES 330, Spring 2020
// 5/2020
// HW 3, Part 1
// Creates a 16 bit counter using T flipflop and
// and gates 
// 412.2 MHz
// The difference between 4 bit counter and 16bit
// counter we CAn have 4 digit number represented 
// in 7 segement display. Also, 16bit counter is 
// combination of 4 4bit counters 
// ISSUES: I have to press Clock 5 times to get from 9 to 10 or 19 to 20 or etc
// Author: Shahzoda Staroverov

module part1(KEY, SW, LEDR, LEDG, HEX0, HEX1, HEX2, HEX3);
	input KEY[0]; //KEY0
	input [1:0] SW; //SW0, SW1
	output [1:0] LEDR; //LEDR0, LEDR 1
	output LEDG[0]; //LEDG0	
	output [6:0] HEX0, HEX1, HEX2, HEX3;// 7 bit vectors for hex values
	assign LEDR = SW; //assign red LEDs to the switch bit 
	assign LEDG[0] = KEY[0]; //assign green LEDs to the switch bit 
	sixteenbitcounter(KEY[0], SW[1], SW[0], HEX0, HEX1, HEX2, HEX3); //calls the module
endmodule 
